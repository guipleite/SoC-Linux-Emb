library IEEE;
use IEEE.std_logic_1164.all;

entity LAB2_FPGA_NIOS is
    port (
        -- Gloabals
        fpga_clk_50        : in  std_logic;             -- clock.clk

        -- I/Os
        fpga_led_pio       : out std_logic_vector(5 downto 0)
  );
end entity LAB2_FPGA_NIOS;

architecture rtl of LAB2_FPGA_NIOS is

component niosLab2 is
  port (
		clk_clk         : in  std_logic                    := 'X'; -- clk
		leds_export     : out std_logic_vector(5 downto 0);        -- export
		reset_reset_n   : in  std_logic                    := 'X'; -- reset_n
		motor_export    : out std_logic_vector(5 downto 0);        -- export
		switches_export : out std_logic_vector(5 downto 0)         -- export
  );
end component niosLab2;

begin


u0 : component niosLab2
  port map (
		clk_clk         => fpga_clk_50,         --      clk.clk
		leds_export     => "!",     --     leds.export
		reset_reset_n   => CONNECTED_TO_reset_reset_n,   --    reset.reset_n
		motor_export    => CONNECTED_TO_motor_export,    --    motor.export
		switches_export => CONNECTED_TO_switches_export  -- switches.export
);


end rtl;


