
module niosLab2 (
	reset_reset_n,
	clk_clk,
	leds_export);	

	input		reset_reset_n;
	input		clk_clk;
	output	[5:0]	leds_export;
endmodule
