
module niosLab2 (
	clk_clk,
	reset_reset_n,
	leds_name);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	leds_name;
endmodule
